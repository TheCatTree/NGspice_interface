*** RF switch circuit ***

* Input source
vs 1 0 dc 0V ac 1V
Rs in 1 50ohm

* Switch
Ci in 4 1.6nF
Rb 4 3 2.1k
Lc1 3 2 100uH
D1 4 5 mydiode
Lc2 5 0 100e-6
cout 5 out 1.6n

* Load
Rload out 0 1000

* DC biasing
vcc 2 0 5V

.model mydiode d (is=1e-15A n=1)

.end